module Ms （）