module test (a,b,c)



endmodule