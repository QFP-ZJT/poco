module module_name (ports)
// 声明
reg,wire,parameter,
input,output,inout,
function,task, ···
// 语句
initial 语句
always  语句
module  实例化
门实例化
用户定义原语(UDP)实例化
连续赋值(Continuous assignment)
endmodule
