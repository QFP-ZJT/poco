/** 
 * ʱ�ӿ���ROM�������������ָ��
 * ��ǰʵ��Ķ������ģ��
 * �̳�ʵ��һ
 */
module test_1(
	input  wire		  in_clk, /*ʱ������Դ*/
	input  wire		  rst,    /*���ָ��  Ϊ0ʱ�����*/
	input  wire 	  run,	  /*�Ƿ�������״̬*/
	input  wire[23:0] in_rom, /*ROM�ڴ����*/
	input  wire[7:0]  keyboard, /*��������*/
	input  wire       interrupt, /*�������� 1��ʱ������*/
	input  wire       in_rom_efficient,/*rom ����ָ����Ч  Ϊ1ʱ��Ч*/
	output wire[7:0]  addr_rom,/*ROM��ַ���*/
	output wire		  out_clk,/*ROM����ָ��*/
	output wire		  wupc,	  /*����ROM���ڶ�״̬*/
	output wire[39:0] led,	  /*led����������*/
    inout  wire[7:0]  dataram, /*����ram*/ 
    output wire[7:0]  addr_ram,/*RAM��ַ���*/
    output wire		  wram,	  /*����RAM����д״̬*/
    output wire		  rram	  /*����ROM���ڶ�״̬*/
);
	/*���߶���*/
	wire [7:0] dbus;		/*CPU�ڲ�����*/

    /*������Ч��romָ������*/
	wire [23:0] in_rom_e;
	wire clk;
    /*�Ĵ���д��������*/
	wire [7:0] reg_ch_w; 	/*д�Ĵ���ѡ����*/
	wire [7:0] reg_ch_r;	/*���Ĵ���ѡ����*/

    /*״̬�Ĵ����������*/
	wire [7:0] reg_sta;		/*״̬������*/

    /*�ۼӼĴ��� �����������*/
	wire [7:0] addtoalu;	/*�ۼ�������ALU*/
	wire [7:0] toans;		/*���ӵ�����Ĵ���*/
	wire [7:0] irtoupc;		/*IR to UPC*/

	//����ʱ���Ƿ�������״̬
	assign clk = run ? in_clk : 1'bz;				/*��runΪtrue �����ʱ�ӣ�����Ͽ�ʱ��*/
	// ROM ����
	assign out_clk = ~clk;						/*cpuIR    �����Ƿ���Ҫȡ��   ����*/
	assign w_uPC = 1'b0;
	assign in_rom_e = in_rom_efficient ? in_rom : 24'b0;
    // RAM ����
    //����ram��dbus
    //assign dbus =  dataram;                     /* ʵ����ȴ���֤������Ƶ���ȷ��  ����̫�����  ����*/
    //ram��ַ����   in_rom_e[5] = 1��ʱ������MAR
    wire [7:0] addr_frommar;
    wire [7:0] addr_frompc;
    // д������
    assign wram = ~in_rom_e[4];
    assign rram = ~in_rom_e[3];

	// ��ʱ�����ʾ
	assign led[7:0] = reg_sta; //(2,2)
	assign led[15:8] = addr_frompc;//(1,2)
	// assign led[23:16] = addr_ram;//�����
	assign led[31:24] = addr_rom;//(1,3)

	// IO ������
	reg [7:0] in_keyboard;
	always@(negedge clk)
	begin
		in_keyboard <= keyboard;
	end
	assign dbus = (in_rom_e[10]==1'b0 && in_rom_e[9] == 1'b1) ? in_keyboard : 8'bz;//IN

	reg [7:0] led_reg;
	assign led[23:16] = led_reg;//(1,1)
	always@(negedge clk)
	begin 
		if(in_rom_e[10]==1'b1 && in_rom_e[9] == 1'b0)
			led_reg <= dbus;
	end


    /*�Ĵ���д��������������*/
    wrcontroller wrcontroller(
        .reg_ch_l   (in_rom_e[15:13]), 	    /*��λָ���ļĴ���ѡ����	(24λ΢�������ָ��)*/
	    .reg_ch_h   (in_rom_e[20:18]), 	    /*��λָ���ļĴ���ѡ����*/
	    .l_wr       (in_rom_e[12:11]),	    /*��λָ���ļĴ��� д��������*/
        .h_wr       (in_rom_e[17:16]),      /*��λָ���ļĴ��� д��������*/
		.next		(in_rom_e[2:0]),		/*����	PCת��	ͣ��*/
	    .reg_ch_w   (reg_ch_w),             /*д�Ĵ���ѡ����*/
	    .reg_ch_r	(reg_ch_r)              /*���Ĵ���ѡ����*/
    );

    /**
     *	ram ��ַ������
     */
     addrforram addrforram(
        .addr_frommar   (addr_frommar),
        .addr_frompc    (addr_frompc),    //ram ��ַ��Դ
        .in_rom_e       (in_rom_e[5]),             //ѡ���ź�
        .addr_ram       (addr_ram)  //��ַ���
     );
	/**
	 * upc��ַ���� 
	 */
	w_uPC upc(
		.clk	(clk),
		.rst	(rst),
		.ld		(in_rom_e[2]),
		.op		(in_rom_e[1:0]),
		.in_upc	(in_rom_e[20:13]),
		.in_pc	(irtoupc),
		.reg_sta(reg_sta),
		.interrupt(interrupt),
		.out	(addr_rom)
	);

	/*
	 *  �Ĵ����ı��
	 *	PC(0) IR(1) MAR(2) MDR(3) ״̬�Ĵ��� �ۼ���(4) ���ݼĴ���(5) ��ַ�Ĵ���(6) R0(7)
	 */
	register reg_add(			/*�ۼӼĴ���*/
		.clk		(clk),
		.in			(dbus),
		.out		(addtoalu),
		.out_allow	(1'b1),
		.in_allow	(reg_ch_w[4]),
		.rst		(rst)
	);

	register reg_ans(			/*�������Ĵ���*/
		.clk		(clk),
		.in			(toans),
		.out		(dbus),
		.out_allow	(reg_ch_r[5]),
		.in_allow	(reg_ch_w[5]),
		.rst		(rst)
	);

	registerformdr reg_mdr(				//ʵ��һ ��ʱ���õ�MDR��ROM��ץȡ����
                                    //ʵ��� mdr��������ԴΪRAM TODO ���� ��ʱȡ��
		.clk		(clk),
		.in			(dbus),
		.out		(dbus),
		.out_allow	(reg_ch_r[3]),		
		.in_allow	(reg_ch_w[3]),
		.ioram		(dataram),
		.rwforram	(in_rom_e[4:3]),
		.rst		(rst),
		.aa			(led[39:32])//(2,3)
	);

    registerforoutput reg_mar(         //MAR�Ĵ���
        .clk		(clk),
		.in			(dbus),
		.inc		(1'b0),
		.out		(dbus),
		.out_allow	(reg_ch_r[2]),		
		.in_allow	(reg_ch_w[2]),
		.rst		(rst),
        .out_direct      (addr_frommar)
    );

    registerforoutput reg_pc(         //PC�Ĵ���
        .clk		(clk),
		.in			(dbus),
		.inc		(in_rom_e[8]),
		.out		(dbus),
		.out_allow	(reg_ch_r[0]),		
		.in_allow	(reg_ch_w[0]),
		.rst		(rst),
        .out_direct      (addr_frompc)
    );

	registerforoutput reg_ir(         //IR�Ĵ���
        .clk		(clk),
		.in			(dbus),
		.inc		(1'b0),
		.out		(dbus),
		.out_allow	(reg_ch_r[1]),		
		.in_allow	(reg_ch_w[1]),
		.rst		(rst),
        .out_direct      (irtoupc)
    );

	register reg_r0(				//ͨ�üĴ���R0
		.clk		(clk),
		.in			(dbus),
		.out		(dbus),
		.out_allow	(reg_ch_r[7]),		
		.in_allow	(reg_ch_w[7]),
		.rst		(rst)
    );

	register reg_r1(				//ͨ�üĴ���R1
		.clk		(clk),
		.in			(dbus),
		.out		(dbus),
		.out_allow	(reg_ch_r[6]),		
		.in_allow	(reg_ch_w[6]),
		.rst		(rst)
	);

    /**
     * alu ���㹦��   ��Ҫ״̬λ�Ľ�Ϊ��־
     */
	w_alu alu(							/*���㵥Ԫ*/
		.clk		(clk),
        .rst        (rst),              /*���*/
		.op			(in_rom_e[23:21]) 	/*ѡ��Ҫִ�еĲ���*/,
		.in_a		(addtoalu)			/*�����ۼ���*/, 
		.in_b		(dbus)				/*����BUS*/,
        .controllerforstate (in_rom_e[7:6]),/*״̬�Ĵ�������λ*/
		.out		(toans)				/*�͵�ans�Ĵ�����*/,
        .mem        (reg_sta)           /*״̬�Ĵ������*/
	);
endmodule



// ΢�������ָ��ĵ�ַ������   
module w_uPC(input clk,input rst,input ld,input [1:0] op,//�µ�ַ���ɷ�ʽ
			input [7:0] reg_sta, 						//״̬�Ĵ���
			input interrupt,							//�ж�
			input [7:0] in_upc,input [7:0] in_pc,output wire [7:0] out);
		/**
		*	rst = 0 ����
		*	rst = 1, ld = 0; ֱ�� out = in
		*		op[1:0] == 01 in_pc;
		*		op[1:0] == 10 in_upc;
		*	rst = 1, ld = 1,op[1:0] == 00; ����
		*	���ܵĸ���:regֱ�����
		*/
		wire [7:0] pctoupc;
		decode_7 decode(
			.in(in_pc),
			.out(pctoupc)
		);
		reg [7:0] value;
		always @(posedge clk) begin
			if (!rst)
				value <= 8'b0;	
			else begin
				case({ld,op[1:0]})	
					3'b100: value <= value + 1;
					3'b001: value <= pctoupc;//����
					3'b010: value <= in_upc; //jump
					3'b000:begin//��������ת
							value <= 8'b0000_0011;
							end
					3'b011: begin//����
							if(reg_sta[2]==1)//�����������  ������������
								value <= 8'b0;
							else
								value <= 8'b0000_0011;		//�������ת��MARָ����λ����
							end
					3'b101: begin
								if(interrupt)
									value <= 8'b0000_0111;
								else
									value <= 8'b0000_0000;
							end
				endcase
			end
		end
		assign out = value;
endmodule


/**
 *	��ͨ�Ĵ������ģ��
 */
module register(
	input clk, input [7:0] in, output wire [7:0] out,
	input out_allow,input in_allow,input rst);

		/** 
		*	rst = 0   ����
		*	in_allow  ��������
		*	out_allow �������
		*/
		reg  [7:0] mem;
		always @(negedge clk) begin
			if (!rst)
				mem <= 8'b00000000;
			else if (in_allow)
				mem <= in;
		end
		assign out = out_allow ? mem : 8'bzzzzzzzz;
endmodule

/** 
 *  MDRר�üĴ��� http://blog.sina.com.cn/s/blog_7bf0c30f0100tedd.html
 */
module registerformdr(
	input clk, input [7:0] in, output wire [7:0] out,
	input out_allow,input in_allow,input rst,
    inout wire [7:0] ioram/*����ram*/,
    input wire [1:0] rwforram /*��ram������ǽ�������*/,
    output wire [7:0] aa
    );

		/** 
		*	rst = 0   ����
		*	in_allow  ��������
		*	out_allow �������
        *   rwforram[1] ioram �������
        *   rwforram[0] ioram ��������
		*/
		reg  [7:0] mem;
		always @(negedge clk) begin
			if (!rst)
				mem <= 8'b0;
			else if (in_allow)
				mem <= in;
			else if (rwforram[0]) //read ram
				mem <= ioram;
		end
		assign out = out_allow ? mem : 8'bzzzzzzzz;

		//д ram
		assign ioram = rwforram[1] ? mem : 8'bz;
		assign aa = mem;
endmodule

/**
 *  for MAR IR PC ר�üĴ���
 */
module registerforoutput(
	input clk, input [7:0] in, input wire inc, output wire [7:0] out,
	input out_allow,input in_allow,input rst, output wire [7:0] out_direct);

		/** 
		*	rst = 0   ����
		*	in_allow  ��������
		*	out_allow �������
		*/
		reg  [7:0] mem;
		always @(negedge clk) begin
			if (!rst)
				mem <= 8'b00000000;
			else if (in_allow)
				mem <= in;
			if(inc)
				mem <= mem+1;
		end
        assign out_direct = mem;
		assign out = out_allow ? mem : 8'bzzzzzzzz;
endmodule

// /**
//  * Ϊ״̬�Ĵ������õ�
//  */
// module registerforstate(
// 	input clk, 
//     input in,
//     input in_allow,
//     output wire [7:0] out,
// 	input rst);

// 		/** 
// 		*	rst = 0   ����
// 		*	in_allow  ��������
// 		*	
// 		*/
		
// endmodule

/**
 * ����߼���ALU��Ƶ�·
 * clk,op ѡ��Ҫִ�еĲ���,
 * in_a�����ۼ���, in_b����BUS,cin��λ��־λ, out���ӵ�����,cout����״̬�Ĵ���
 */
module w_alu (
	input clk, input rst,input [2:0] op/*ѡ��Ҫִ�еĲ���*/,input [7:0] in_a/*�����ۼ���*/, input [7:0] in_b/*����BUS*/,
    input wire [1:0] controllerforstate,/*״̬�Ĵ���������*/
	output reg [7:0] out/*���ӵ�����*/,output reg [7:0] mem/*״̬�Ĵ��������*/);
		/**
		*	op 000 �ӷ�
		*	op 001 ����
		*	op 010 �˷�
		*	op 011 ��in_bȡ��	
		*	op 100 in_a,in_b���
		*	op 101 in_b,����1     ΪPC����
		*	op 110 ����
		*	op 111 �����
        *
        *   ״̬�Ĵ��� �����ȫΪ0 ���ж����յĽ����Ϊ1   �����
		*/
        wire [7:0] in_allow;
        reg cout_add;reg cout_sub;
        wire equal;/*�ж�����Ƿ�Ϊȫ0*/
        assign equal = out[0] | out[1] | out[2] | out[3] | out[4] | out[5] | out[6] | out[7];
			   /** ״̬λ����
				* 0:	��λ��־�� 
				* 1:	��λ��־��
				* 2:	���Ϊ0 Ϊ1
				* 3:   �������������
				* 4:   �������㸺���
				*/
		always @(*) begin
            if (!rst)
				mem <= 8'b0;
			case(op)//ʹ��˫����λ�Ĳ����������
				3'b000:	begin       //�ӷ�
				 	case(controllerforstate)
					2'b00:begin
						{cout_add,out[7:0]} <= {in_a[7],in_a}+{in_b[7],in_b};
						if({cout_add,out[7]} == 2'b01) // ����
							mem[3] <= 1'b1;
						if({cout_add,out[7]} == 2'b10) //����
							mem[4] <= 1'b1;
						end
					2'b01:{mem[0],out[7:0]} <= {in_a}+{in_b};//��¼��λ
					2'b10:begin out[7:0] <= {in_a}+{in_b};//ʹ�ý�λ
							   out[7:0] <= out[7:0] + mem[0];
						 end
					2'b11:{mem[0],out[7:0]} <= {in_a}+{in_b}+{7'b0000000,mem[0]};//��¼��ʹ�ý�λ
					endcase
					mem[2] <= ~equal;
					end
				3'b001:  begin       //����
						{cout_sub,out[7:0]} <= {in_a[7],in_a}+{~in_b[7],~in_b}+9'd1;
						if({cout_add,out[7]} == 2'b01) // ����
							mem[3] <= 1'b1;
						if({cout_add,out[7]} == 2'b10) //����
							mem[4] <= 1'b1;
						mem[2] <= ~equal;
					end
				3'b010:  begin out[7:0] <= in_a*in_b;mem[2] <= ~equal;end
				3'b011:  begin out[7:0] <= ~in_b;mem[2] <= ~equal;end
				3'b100:  begin out[7:0] <= in_a^in_b;mem[2] <= ~equal;end
				3'b101:  begin out[7:0] <= in_b+1;mem[2] <= ~equal;end
                3'b110:  begin out[7:0] <= in_a / in_b;mem[2] <= ~equal;end
				3'b111:  out[7:0] <= 8'bz;
			endcase	
			
		end
endmodule


/**
 * RAM ��ַ���
 */
module addrforram(
    input [7:0] addr_frommar,
    input [7:0] addr_frompc,    //ram ��ַ��Դ
    input in_rom_e,             //ѡ���ź�
    output wire [7:0] addr_ram  //��ַ���
    );
    assign addr_ram = in_rom_e ? addr_frommar : addr_frompc;
endmodule



/**
 *  �Ĵ���д��������    ������߼�
 */
module wrcontroller(
    input [2:0] reg_ch_l, 	    /*��λָ���ļĴ���ѡ����	(24λ΢�������ָ��)*/
	input [2:0] reg_ch_h, 	    /*��λָ���ļĴ���ѡ����*/
	input [1:0] l_wr,	        /*��λָ���ļĴ��� д��������*/
    input [1:0] h_wr,           /*��λָ���ļĴ��� д��������*/
	input [2:0] next,		    /*�����µ�ַ���ɷ�ʽ�����Ƿ���Ч*/
	output wire [7:0] reg_ch_w, /*д�Ĵ���ѡ����*/
	output wire [7:0] reg_ch_r	/*���Ĵ���ѡ����*/);

    wire [7:0] reg_ch_l_w; 	/*��λָ����д�Ĵ���ѡ����	(24λ΢�������ָ��)*/
	wire [7:0] reg_ch_l_r;	/*��λָ���Ķ��Ĵ���ѡ����*/
	wire [7:0] reg_ch_h_w; 	/*��λָ����д�Ĵ���ѡ����*/
	wire [7:0] reg_ch_h_r;	/*��λָ���Ķ��Ĵ���ѡ����*/

    decode decode_l_r(			/*��λָ���Ķ��Ĵ���*/
		.in 	(reg_ch_l),
		.open	(l_wr[0]),
		.out 	(reg_ch_l_r)
	);
	decode decode_l_w(			/*��λָ����д�Ĵ���*/
		.in 	(reg_ch_l),
		.open	(l_wr[1]),
		.out 	(reg_ch_l_w)
	);
	decode decode_2_r(			/*��λָ���Ķ��Ĵ���*/
		.in 	(reg_ch_h),
		.open	(h_wr[0]),
		.out 	(reg_ch_h_r)
	);
	decode decode_2_w(			/*��λָ����д�Ĵ���*/
		.in 	(reg_ch_h),
		.open	(h_wr[1]),
		.out 	(reg_ch_h_w)
	);
    // �Ĵ���״̬������
	//                           ����        ͨ��PCת��        ͣ��
	assign reg_ch_w = (next == 3'b100 || next == 3'b001 || 3'b111) ? (reg_ch_l_w | reg_ch_h_w) : 8'b0; /*д�߻���*/
	assign reg_ch_r = (next == 3'b100 || next == 3'b001 || 3'b111) ? (reg_ch_l_r | reg_ch_h_r) : 8'b0;  /*���߻���*/

endmodule

/**
 *	������  �� - ��   ���ҽ���openΪ1��ʱ��
 */
module decode(
	input [2:0] in,
	input open,
	output reg [7:0] out);
	always @(*)
		if (open)
			case(in)
			3'b000:  out <= 8'b00000001;
			3'b001:  out <= 8'b00000010;
			3'b010:  out <= 8'b00000100;
			3'b011:  out <= 8'b00001000;
			3'b100:  out <= 8'b00010000;
			3'b101:  out <= 8'b00100000;
			3'b110:  out <= 8'b01000000;
			3'b111:  out <= 8'b10000000;
			endcase
		else
			out <= 8'b00000000;
endmodule

/**
 *
 */
module decode_7(
	input [7:0] in,
	output reg [7:0] out);
	always @(*)
		case(in)
		8'b00110111: out <= 8'b10001010;	// 00110111 TO 138 	ALU_��_R1
8'b00010111: out <= 8'b01010001;	// 00010111 TO 81 	STORE_PC_ANS
8'b00110110: out <= 8'b01111100;	// 00110110 TO 124 	ALU_��_R0
8'b00010000: out <= 8'b00110110;	// 00010000 TO 54 	STORE_MAR_R0
8'b00010010: out <= 8'b00111100;	// 00010010 TO 60 	STORE_MAR_MAR
8'b00010001: out <= 8'b00111001;	// 00010001 TO 57 	STORE_MAR_R1
8'b00100111: out <= 8'b01101100;	// 00100111 TO 108 	R1--PC
8'b00100101: out <= 8'b01101000;	// 00100101 TO 104 	R1--LJ
8'b00001001: out <= 8'b00101101;	// 00001001 TO 45 	LOAD_NUM_R1
8'b00010110: out <= 8'b01001100;	// 00010110 TO 76 	STORE_PC_MAR
8'b00001000: out <= 8'b00101010;	// 00001000 TO 42 	LOAD_NUM_R0
8'b01100001: out <= 8'b10011101;	// 01100001 TO 157 	ALU_��RU_R0
8'b00110101: out <= 8'b10001000;	// 00110101 TO 136 	ALU_��_R1
8'b01100000: out <= 8'b10010111;	// 01100000 TO 151 	ALU_��RU_R1
8'b00110100: out <= 8'b01111010;	// 00110100 TO 122 	ALU_��_R0
8'b01000001: out <= 8'b10011001;	// 01000001 TO 153 	ALU_��R_R0
8'b01000000: out <= 8'b10010011;	// 01000000 TO 147 	ALU_��R_R1
8'b00100011: out <= 8'b01100100;	// 00100011 TO 100 	R0--PC
8'b00100001: out <= 8'b01100000;	// 00100001 TO 96 	R0--LJ
8'b00011000: out <= 8'b01010110;	// 00011000 TO 86 	STORE_NUM_MAR
8'b00100000: out <= 8'b01011110;	// 00100000 TO 94 	RO--MAR
8'b00101000: out <= 8'b01101110;	// 00101000 TO 110 	ANS--MAR
8'b00111010: out <= 8'b10000000;	// 00111010 TO 128 	ALU_����_R0
8'b00111011: out <= 8'b10001110;	// 00111011 TO 142 	ALU_����_R1
8'b10000000: out <= 8'b00000000;	// 10000000 TO 0 	GETPC
8'b00100010: out <= 8'b01100010;	// 00100010 TO 98 	RO--R1
8'b01110110: out <= 8'b10100101;	// 01110110 TO 165 	IN_MAR
8'b00101001: out <= 8'b01110000;	// 00101001 TO 112 	ANS--R1
8'b00000101: out <= 8'b00011011;	// 00000101 TO 27 	LOAD_PC_R1
8'b00101010: out <= 8'b01110010;	// 00101010 TO 114 	ANS--R0
8'b01010000: out <= 8'b10010101;	// 01010000 TO 149 	ALU_��U_R1
8'b00000100: out <= 8'b00010110;	// 00000100 TO 22 	LOAD_PC_R0
8'b00100100: out <= 8'b01100110;	// 00100100 TO 102 	R1--MAR
8'b01010001: out <= 8'b10011011;	// 01010001 TO 155 	ALU_��U_R0
8'b00111000: out <= 8'b01111110;	// 00111000 TO 126 	ALU_���_R0
8'b00111001: out <= 8'b10001100;	// 00111001 TO 140 	ALU_���_R1
8'b00001011: out <= 8'b00110011;	// 00001011 TO 51 	LOAD_NUM_MAR
8'b00010101: out <= 8'b01000111;	// 00010101 TO 71 	STORE_PC_R1
8'b00010100: out <= 8'b01000010;	// 00010100 TO 66 	STORE_PC_R0
8'b00111101: out <= 8'b10010000;	// 00111101 TO 144 	ALU_��_R1
8'b00111100: out <= 8'b10000010;	// 00111100 TO 130 	ALU_��_R0
8'b01111011: out <= 8'b10101011;	// 01111011 TO 171 	OUT_MAR
8'b10000010: out <= 8'b00000111;	// 10000010 TO 7 	CH_INTERRUPT
8'b01110101: out <= 8'b10100001;	// 01110101 TO 161 	IN_R1
8'b01110100: out <= 8'b10011111;	// 01110100 TO 159 	IN_R0
8'b01111010: out <= 8'b10101101;	// 01111010 TO 173 	OUT_ANS
8'b00000110: out <= 8'b00100000;	// 00000110 TO 32 	LOAD_PC_LJ
8'b10000001: out <= 8'b00000011;	// 10000001 TO 3 	GETMAR
8'b11110000: out <= 8'b10010010;	// 11110000 TO 146 	ͣ��
8'b00000010: out <= 8'b00010000;	// 00000010 TO 16 	LOAD_MAR_LJ
8'b00110011: out <= 8'b10000110;	// 00110011 TO 134 	ALU_��_R1
8'b00110010: out <= 8'b01111000;	// 00110010 TO 120 	ALU_��_R0
8'b00000111: out <= 8'b00100101;	// 00000111 TO 37 	LOAD_PC_MAR
8'b10000100: out <= 8'b00001001;	// 10000100 TO 9 	JUMP_N
8'b00100110: out <= 8'b01101010;	// 00100110 TO 106 	R1--R0
8'b00000011: out <= 8'b00010011;	// 00000011 TO 19 	LOAD_MAR_MAR
8'b00001010: out <= 8'b00110000;	// 00001010 TO 48 	LOAD_NUM_LJ
8'b01111000: out <= 8'b10100111;	// 01111000 TO 167 	OUT_R0
8'b10000011: out <= 8'b00001000;	// 10000011 TO 8 	JUMP_E
8'b00011001: out <= 8'b01011001;	// 00011001 TO 89 	STORE_NUM_PC
8'b00101011: out <= 8'b01110100;	// 00101011 TO 116 	ANS--PC
8'b00110001: out <= 8'b10000100;	// 00110001 TO 132 	ALU_��_R1
8'b00110000: out <= 8'b01110110;	// 00110000 TO 118 	ALU_��_R0
8'b01110111: out <= 8'b10100011;	// 01110111 TO 163 	IN_LJ
8'b01111001: out <= 8'b10101001;	// 01111001 TO 169 	OUT_R1
8'b00000000: out <= 8'b00001010;	// 00000000 TO 10 	LOAD_MAR_R0
8'b00000001: out <= 8'b00001101;	// 00000001 TO 13 	LOAD_MAR_R1
8'b00010011: out <= 8'b00111111;	// 00010011 TO 63 	STORE_MAR_ANS
		endcase
endmodule